//
//
// $Id: fw_tb4.v,v 1.1 2005/10/03 21:01:33 osc0414 Exp $
//
// FW Test bench 32x32 matrix
//
// Tests functionality under real conditions for a 32x32 matrix
// Pipeline bubbles 
//
// Uday Kumar Reddy Bondhugula
//
//
//

module fw_tb4;

reg reset;
wire clk;

reg [63:0] fw_in;
reg in_valid;
reg [1:0] phase;

clock   clock(.reset(reset), .clk(clk));

fw		fw_inst(
	.reset(reset),
	.clk(clk),
	.phase(phase),
	.inhibit(),

	.inD(fw_in),
	.in_valid(in_valid),

	.outD(),
	.out_valid()
);

initial
begin
	reset = 1;
	in_valid = 0;
	phase = 2'b00;
	#10 reset = 0;
	#30 reset = 1;
	#10 reset = 0;
end

initial
begin: fw_input
	#65 in_valid = 1;

	// Input an 32x32 matrix
	//
	fw_in =     64'h004e_0057_0054_0000;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 1;
	fw_in = 64'h0057_0024_005e_0010;
	#10 fw_in = 64'h003f_0016_0032_005d;
	#10 fw_in = 64'h0040_003c_005b_001c;
	#10 fw_in = 64'h0049_001b_0029_001b;
	#10 fw_in = 64'h0044_0045_000c_0025;
	#10 fw_in = 64'h003f_001f_0053_001e;
	#10 fw_in = 64'h001e_0024_0044_0018;


	#10 fw_in = 64'h0045_0055_0003_0000;
	#10 fw_in = 64'h002c_004b_002e_0062;
	#10 fw_in = 64'h0019_0058_0020_000c;
	#10 fw_in = 64'h0034_0035_0009_0050;
	#10 fw_in = 64'h003c_0058_005f_002a;
	#10 fw_in = 64'h001d_0017_0005_004b;
	#10 fw_in = 64'h0019_0042_001f_0044;
	#10 fw_in = 64'h004d_0053_0058_0052;


	#10 fw_in = 64'h003b_0017_0000_0003;
	#10 fw_in = 64'h0039_005e_0044_0046;
	#10 fw_in = 64'h004a_001e_002b_000c;
	#10 fw_in = 64'h0026_0055_0014_0016;
	#10 fw_in = 64'h0047_0010_0019_0063;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 1;
	fw_in = 64'h0051_005c_001b_000e;
	#10 fw_in = 64'h0047_003f_004a_0039;
	#10 fw_in = 64'h001a_0006_0052_0061;


	#10 fw_in = 64'h0028_001c_0000_0054;
	#10 fw_in = 64'h0047_0016_002f_0048;
	#10 fw_in = 64'h0017_000d_0052_000b;
	#10 fw_in = 64'h0024_0061_003b_0046;
	#10 fw_in = 64'h0013_0059_0011_0046;
	#10 fw_in = 64'h001a_0053_004d_005c;
	#10 fw_in = 64'h000a_0030_004a_001b;
	#10 fw_in = 64'h0064_0016_0021_0004;


	#10 fw_in = 64'h0025_0000_001c_0055;
	#10 fw_in = 64'h000e_001e_002f_0006;
	#10 fw_in = 64'h0053_0060_0019_003a;
	#10 fw_in = 64'h0023_0044_000f_002e;
	#10 fw_in = 64'h0058_0033_002c_0041;
	#10 fw_in = 64'h0059_004f_004d_0009;
	#10 fw_in = 64'h0037_0034_0004_0055;
	#10 fw_in = 64'h004d_003d_0021_0064;


	#10 fw_in = 64'h000d_0000_0017_0057;
	#10 fw_in = 64'h0054_003b_0034_0052;
	#10 fw_in = 64'h0046_0031_001f_0006;
	#10 fw_in = 64'h0023_004c_0063_004a;
	#10 fw_in = 64'h0027_0027_0035_001b;
	#10 fw_in = 64'h005c_0012_0054_0030;
	#10 fw_in = 64'h0028_0048_000f_0040;
	#10 fw_in = 64'h0035_000b_0053_0015;


	#10 fw_in = 64'h0000_000d_0028_0045;
	#10 fw_in = 64'h0028_005f_0057_001b;
	#10 fw_in = 64'h004f_0023_0047_0060;
	#10 fw_in = 64'h0003_0062_0002_0044;
	#10 fw_in = 64'h0039_0035_005d_0012;
	#10 fw_in = 64'h002a_0057_0051_0002;
	#10 fw_in = 64'h0014_002d_005a_0042;
	#10 fw_in = 64'h0012_0020_001e_0029;


	#10 fw_in = 64'h0000_0025_003b_004e;
	#10 fw_in = 64'h005b_0060_0016_004c;
	#10 fw_in = 64'h0061_0049_0022_0002;
	#10 fw_in = 64'h0028_0059_0025_004d;
	#10 fw_in = 64'h001a_0043_004f_0021;
	#10 fw_in = 64'h000b_001f_0008_0034;
	#10 fw_in = 64'h0001_004d_003c_004e;
	#10 fw_in = 64'h0020_0038_0016_0022;


	#10 fw_in = 64'h004c_0052_0048_0062;
	#10 fw_in = 64'h0044_001c_000a_0000;
	#10 fw_in = 64'h0057_0036_0062_0039;
	#10 fw_in = 64'h0014_0054_0007_0042;
	#10 fw_in = 64'h0021_0048_001d_0019;
	#10 fw_in = 64'h0047_0014_0004_001e;
	#10 fw_in = 64'h0029_0010_0009_0045;
	#10 fw_in = 64'h0013_0018_0061_0032;


	#10 fw_in = 64'h001b_0006_0046_0010;
	#10 fw_in = 64'h0064_001e_0038_0000;
	#10 fw_in = 64'h0052_003c_005f_003e;
	#10 fw_in = 64'h005d_003a_0009_0033;
	#10 fw_in = 64'h0059_0047_001e_003e;
	#10 fw_in = 64'h0013_005e_003c_0020;
	#10 fw_in = 64'h004f_0046_0017_0061;
	#10 fw_in = 64'h0058_0059_0043_0053;


	#10 fw_in = 64'h0016_0034_002f_002e;
	#10 fw_in = 64'h0059_0050_0000_0038;
	#10 fw_in = 64'h0033_002a_001d_0041;
	#10 fw_in = 64'h0041_0023_0001_005e;
	#10 fw_in = 64'h0039_0058_000f_0019;
	#10 fw_in = 64'h0042_001c_005c_002c;
	#10 fw_in = 64'h0034_0021_0025_003c;
	#10 fw_in = 64'h0008_004c_001d_0026;


	#10 fw_in = 64'h0057_002f_0044_005e;
	#10 fw_in = 64'h0049_0026_0000_000a;
	#10 fw_in = 64'h001f_000a_003d_001f;
	#10 fw_in = 64'h0010_001e_0036_0038;
	#10 fw_in = 64'h004b_0055_002f_002b;
	#10 fw_in = 64'h0012_004b_003a_0016;
	#10 fw_in = 64'h000a_0013_0030_0052;
	#10 fw_in = 64'h004e_001a_0040_0052;


	#10 fw_in = 64'h0060_003b_0016_004b;
	#10 fw_in = 64'h0024_0000_0026_001e;
	#10 fw_in = 64'h002c_001d_0013_005e;
	#10 fw_in = 64'h004d_001e_001d_000c;
	#10 fw_in = 64'h000e_0040_002c_0005;
	#10 fw_in = 64'h0005_0029_0007_0027;
	#10 fw_in = 64'h0046_0059_001d_0013;
	#10 fw_in = 64'h0019_0061_0012_0012;


	#10 fw_in = 64'h005f_001e_005e_0024;
	#10 fw_in = 64'h001a_0000_0050_001c;
	#10 fw_in = 64'h0055_0025_0040_004f;
	#10 fw_in = 64'h001c_0025_0031_003d;
	#10 fw_in = 64'h0022_0039_005b_003d;
	#10 fw_in = 64'h0025_001b_002d_0026;
	#10 fw_in = 64'h0036_0002_0019_0042;
	#10 fw_in = 64'h0064_0010_003d_0058;


	#10 fw_in = 64'h005b_0054_0047_002c;
	#10 fw_in = 64'h0000_001a_0049_0064;
	#10 fw_in = 64'h0028_0006_005b_002d;
	#10 fw_in = 64'h0053_0046_0057_0037;
	#10 fw_in = 64'h0008_0062_0041_002b;
	#10 fw_in = 64'h000c_0031_0005_0038;
	#10 fw_in = 64'h002c_0064_001d_0017;
	#10 fw_in = 64'h0017_0029_0045_002f;


	#10 fw_in = 64'h0028_000e_0039_0057;
	#10 fw_in = 64'h0000_0024_0059_0044;
	#10 fw_in = 64'h005d_000b_0064_0006;
	#10 fw_in = 64'h0005_003d_0004_002b;
	#10 fw_in = 64'h003a_0012_0030_0012;
	#10 fw_in = 64'h0040_005e_0064_0029;
	#10 fw_in = 64'h0052_0004_0053_003d;
	#10 fw_in = 64'h003a_0047_0053_0010;


	#10 fw_in = 64'h0002_0006_000b_000c;
	#10 fw_in = 64'h0006_004f_001f_003e;
	#10 fw_in = 64'h002d_0025_0015_0000;
	#10 fw_in = 64'h0009_0042_0017_001b;
	#10 fw_in = 64'h0019_003b_0053_0011;
	#10 fw_in = 64'h0001_0019_003f_0026;
	#10 fw_in = 64'h0050_0064_0035_0025;
	#10 fw_in = 64'h004a_0048_0045_0033;


	#10 fw_in = 64'h0060_003a_000c_005d;
	#10 fw_in = 64'h002d_005e_0041_0039;
	#10 fw_in = 64'h0049_002b_0052_0000;
	#10 fw_in = 64'h001e_000f_0022_0050;
	#10 fw_in = 64'h0052_0007_0047_0018;
	#10 fw_in = 64'h0038_0057_000c_0037;
	#10 fw_in = 64'h000f_0036_0024_0025;
	#10 fw_in = 64'h0043_0026_000c_0061;


	#10 fw_in = 64'h0022_001f_0052_0020;
	#10 fw_in = 64'h0064_0040_003d_005f;
	#10 fw_in = 64'h0061_0064_0000_0052;
	#10 fw_in = 64'h0045_000e_004a_003c;
	#10 fw_in = 64'h0043_001b_0060_005b;
	#10 fw_in = 64'h0055_005b_0029_0055;
	#10 fw_in = 64'h0008_0025_002b_004d;
	#10 fw_in = 64'h0013_0050_0039_002e;


	#10 fw_in = 64'h0047_0019_002b_0032;
	#10 fw_in = 64'h005b_0013_001d_0062;
	#10 fw_in = 64'h0049_0058_0000_0015;
	#10 fw_in = 64'h0032_0016_0022_0055;
	#10 fw_in = 64'h005e_003d_0034_003e;
	#10 fw_in = 64'h005b_0036_001c_001f;
	#10 fw_in = 64'h0027_0022_0021_0038;
	#10 fw_in = 64'h0035_0036_0056_001a;


	#10 fw_in = 64'h0049_0031_000d_0058;
	#10 fw_in = 64'h000b_0025_000a_003c;
	#10 fw_in = 64'h0007_0000_0058_002b;
	#10 fw_in = 64'h0016_0049_000e_0002;
	#10 fw_in = 64'h0016_0064_0014_0038;
	#10 fw_in = 64'h0029_000c_0028_0005;
	#10 fw_in = 64'h001c_001d_0006_0044;
	#10 fw_in = 64'h0015_003b_0055_0033;


	#10 fw_in = 64'h0023_0060_001e_0016;
	#10 fw_in = 64'h0006_001d_002a_0036;
	#10 fw_in = 64'h0033_0000_0064_0025;
	#10 fw_in = 64'h0041_003d_0031_005e;
	#10 fw_in = 64'h003b_0032_0051_0052;
	#10 fw_in = 64'h003b_002c_0033_0063;
	#10 fw_in = 64'h005a_0008_0005_0047;
	#10 fw_in = 64'h0012_0009_0057_0005;


	#10 fw_in = 64'h0061_0046_0017_0019;
	#10 fw_in = 64'h005d_0055_001f_0052;
	#10 fw_in = 64'h0000_0033_0049_0049;
	#10 fw_in = 64'h0064_0017_0056_001a;
	#10 fw_in = 64'h000e_0063_002b_0029;
	#10 fw_in = 64'h005b_0019_005b_0063;
	#10 fw_in = 64'h0025_0014_0052_000a;
	#10 fw_in = 64'h0005_005f_0038_0021;


	#10 fw_in = 64'h004f_0053_004a_003f;
	#10 fw_in = 64'h0028_002c_0033_0057;
	#10 fw_in = 64'h0000_0007_0061_002d;
	#10 fw_in = 64'h0056_0005_005b_0006;
	#10 fw_in = 64'h0047_0026_0020_000a;
	#10 fw_in = 64'h001f_004b_0025_001a;
	#10 fw_in = 64'h001b_003c_0037_0013;
	#10 fw_in = 64'h002a_0017_0056_0017;


	#10 fw_in = 64'h004d_004a_0046_0050;
	#10 fw_in = 64'h002b_003d_0038_0033;
	#10 fw_in = 64'h0006_005e_0055_0050;
	#10 fw_in = 64'h0005_0044_0016_0000;
	#10 fw_in = 64'h001b_0037_003e_000e;
	#10 fw_in = 64'h0003_0003_002d_003c;
	#10 fw_in = 64'h002b_0016_0055_0007;
	#10 fw_in = 64'h0049_005a_001d_0045;


	#10 fw_in = 64'h0044_002e_0016_001c;
	#10 fw_in = 64'h0037_000c_005e_0042;
	#10 fw_in = 64'h001a_0002_003c_001b;
	#10 fw_in = 64'h001e_001d_0037_0000;
	#10 fw_in = 64'h0064_0006_005e_005b;
	#10 fw_in = 64'h0005_000f_003d_0052;
	#10 fw_in = 64'h0044_001d_002c_000c;
	#10 fw_in = 64'h0024_0054_001f_005d;


	#10 fw_in = 64'h0025_0063_003b_0009;
	#10 fw_in = 64'h0004_0031_0036_0009;
	#10 fw_in = 64'h005b_0031_0022_0022;
	#10 fw_in = 64'h002f_0044_0000_0037;
	#10 fw_in = 64'h002f_0001_001e_0045;
	#10 fw_in = 64'h005b_0032_0062_0059;
	#10 fw_in = 64'h0062_0040_0022_0004;
	#10 fw_in = 64'h001a_0057_005d_0036;


	#10 fw_in = 64'h0002_000f_0014_005b;
	#10 fw_in = 64'h0057_001d_0001_0007;
	#10 fw_in = 64'h0056_000e_004a_0017;
	#10 fw_in = 64'h002c_001c_0000_0016;
	#10 fw_in = 64'h0012_003c_003a_001a;
	#10 fw_in = 64'h0048_000e_0013_0011;
	#10 fw_in = 64'h0030_0007_0063_002b;
	#10 fw_in = 64'h0045_0033_005b_0034;


	#10 fw_in = 64'h0059_004c_0061_0035;
	#10 fw_in = 64'h003d_0025_001e_003a;
	#10 fw_in = 64'h0005_003d_0016_000f;
	#10 fw_in = 64'h0033_0000_001c_001d;
	#10 fw_in = 64'h005f_0003_0039_0031;
	#10 fw_in = 64'h0028_002c_0064_0062;
	#10 fw_in = 64'h0001_0004_001d_0003;
	#10 fw_in = 64'h003c_0027_0030_0052;


	#10 fw_in = 64'h0062_0044_0055_003c;
	#10 fw_in = 64'h0046_001e_0023_0054;
	#10 fw_in = 64'h0017_0049_000e_0042;
	#10 fw_in = 64'h0024_0000_0044_0044;
	#10 fw_in = 64'h0028_0012_001c_0061;
	#10 fw_in = 64'h003e_0050_0006_0011;
	#10 fw_in = 64'h0018_0062_0057_0021;
	#10 fw_in = 64'h0063_003a_0054_0062;


	#10 fw_in = 64'h0028_0023_0024_0034;
	#10 fw_in = 64'h0005_001c_0010_005d;
	#10 fw_in = 64'h0056_0041_0032_001e;
	#10 fw_in = 64'h0000_0024_002c_001e;
	#10 fw_in = 64'h0048_0027_0001_004e;
	#10 fw_in = 64'h0059_0044_005a_0032;
	#10 fw_in = 64'h002d_002c_0060_005d;
	#10 fw_in = 64'h0029_0053_005b_001e;


	#10 fw_in = 64'h0003_0023_0026_0040;
	#10 fw_in = 64'h0053_004d_0041_0014;
	#10 fw_in = 64'h0064_0016_0045_0009;
	#10 fw_in = 64'h0000_0033_002f_0005;
	#10 fw_in = 64'h0046_0013_000d_0044;
	#10 fw_in = 64'h0022_004e_0040_0003;
	#10 fw_in = 64'h0058_0015_0029_0061;
	#10 fw_in = 64'h0055_0062_000f_0021;


	#10 fw_in = 64'h0021_001b_0046_002a;
	#10 fw_in = 64'h0012_003d_002b_003e;
	#10 fw_in = 64'h000a_0052_003e_0018;
	#10 fw_in = 64'h0044_0061_001a_005b;
	#10 fw_in = 64'h005b_0023_004e_0000;
	#10 fw_in = 64'h000f_003a_0019_001b;
	#10 fw_in = 64'h000d_003b_0006_0045;
	#10 fw_in = 64'h001b_002f_0001_0057;


	#10 fw_in = 64'h0012_0041_0063_001b;
	#10 fw_in = 64'h002b_0005_0019_0019;
	#10 fw_in = 64'h0029_0038_005b_0011;
	#10 fw_in = 64'h004e_0031_0045_000e;
	#10 fw_in = 64'h0040_002e_0057_0000;
	#10 fw_in = 64'h0056_003f_0032_0020;
	#10 fw_in = 64'h0020_0055_004f_0050;
	#10 fw_in = 64'h0060_001c_004d_0023;


	#10 fw_in = 64'h004f_0035_0011_005f;
	#10 fw_in = 64'h0030_005b_002f_001e;
	#10 fw_in = 64'h0020_0051_0034_0047;
	#10 fw_in = 64'h000d_001c_003a_005e;
	#10 fw_in = 64'h0038_000f_0000_0057;
	#10 fw_in = 64'h0050_000d_005b_000d;
	#10 fw_in = 64'h004b_005a_0046_000b;
	#10 fw_in = 64'h0022_0015_002a_0038;


	#10 fw_in = 64'h005d_002c_0019_0029;
	#10 fw_in = 64'h0041_002c_000f_001d;
	#10 fw_in = 64'h002b_0014_0060_0053;
	#10 fw_in = 64'h0001_0039_001e_003e;
	#10 fw_in = 64'h0017_0054_0000_004e;
	#10 fw_in = 64'h005a_004c_002d_0028;
	#10 fw_in = 64'h0021_0009_003c_0016;
	#10 fw_in = 64'h004d_001b_0011_0052;


	#10 fw_in = 64'h0043_0027_0059_0058;
	#10 fw_in = 64'h0012_0039_0055_0047;
	#10 fw_in = 64'h0026_0032_003d_0007;
	#10 fw_in = 64'h0013_0012_003c_0006;
	#10 fw_in = 64'h004a_0000_0054_002e;
	#10 fw_in = 64'h005a_0026_004a_003b;
	#10 fw_in = 64'h003a_004f_0008_0054;
	#10 fw_in = 64'h0001_001e_0048_000f;


	#10 fw_in = 64'h0035_0033_0010_001b;
	#10 fw_in = 64'h0062_0040_0058_0048;
	#10 fw_in = 64'h0063_0064_001b_003b;
	#10 fw_in = 64'h0027_0003_0001_0037;
	#10 fw_in = 64'h005f_0000_000f_0023;
	#10 fw_in = 64'h004a_0059_000c_0061;
	#10 fw_in = 64'h0017_0023_003f_0047;
	#10 fw_in = 64'h0006_0046_0015_0007;


	#10 fw_in = 64'h001a_0027_0013_003c;
	#10 fw_in = 64'h003a_0022_004b_0059;
	#10 fw_in = 64'h0047_003b_005e_0052;
	#10 fw_in = 64'h0046_0028_0012_0064;
	#10 fw_in = 64'h0000_005f_0017_0040;
	#10 fw_in = 64'h003f_0020_0030_004a;
	#10 fw_in = 64'h005c_005d_005b_0053;
	#10 fw_in = 64'h003a_0016_0010_003a;


	#10 fw_in = 64'h0039_0058_0047_0049;
	#10 fw_in = 64'h0008_000e_0039_0021;
	#10 fw_in = 64'h000e_0016_0043_0019;
	#10 fw_in = 64'h0048_005f_002f_001b;
	#10 fw_in = 64'h0000_004a_0038_005b;
	#10 fw_in = 64'h0005_0014_0006_0005;
	#10 fw_in = 64'h0052_0063_003f_0055;
	#10 fw_in = 64'h0043_0048_005d_0010;


	#10 fw_in = 64'h0034_0030_005c_004b;
	#10 fw_in = 64'h0029_0026_0016_0020;
	#10 fw_in = 64'h001a_0063_001f_0037;
	#10 fw_in = 64'h0003_0011_0011_0052;
	#10 fw_in = 64'h0005_0061_0028_0020;
	#10 fw_in = 64'h0013_0051_0027_0000;
	#10 fw_in = 64'h000d_003f_0047_0016;
	#10 fw_in = 64'h0025_0056_004e_0050;


	#10 fw_in = 64'h0002_0009_000e_0025;
	#10 fw_in = 64'h0038_0027_002c_001e;
	#10 fw_in = 64'h0063_0005_0055_0026;
	#10 fw_in = 64'h0032_0062_0059_003c;
	#10 fw_in = 64'h004a_003b_000d_001b;
	#10 fw_in = 64'h0034_000b_0023_0000;
	#10 fw_in = 64'h004c_005c_0054_0049;
	#10 fw_in = 64'h001d_0034_001a_003a;


	#10 fw_in = 64'h0008_0054_004d_0005;
	#10 fw_in = 64'h0064_002d_003a_003c;
	#10 fw_in = 64'h0025_0033_001c_000c;
	#10 fw_in = 64'h0040_0006_0013_003d;
	#10 fw_in = 64'h0006_000c_002d_0032;
	#10 fw_in = 64'h004c_005c_0000_0023;
	#10 fw_in = 64'h0045_005a_000f_0038;
	#10 fw_in = 64'h0053_0006_0013_005e;


	#10 fw_in = 64'h0051_004d_001b_000c;
	#10 fw_in = 64'h0005_0007_005c_0004;
	#10 fw_in = 64'h005b_0028_0029_003f;
	#10 fw_in = 64'h005a_0064_0062_002d;
	#10 fw_in = 64'h0030_004a_005b_0019;
	#10 fw_in = 64'h0006_0021_0000_0027;
	#10 fw_in = 64'h0033_004d_002a_001c;
	#10 fw_in = 64'h0037_0032_001d_0009;


	#10 fw_in = 64'h001f_0012_0053_0017;
	#10 fw_in = 64'h005e_001b_004b_005e;
	#10 fw_in = 64'h004b_002c_0036_0057;
	#10 fw_in = 64'h004e_0050_000e_000f;
	#10 fw_in = 64'h0014_0059_004c_003f;
	#10 fw_in = 64'h005f_0000_0021_000b;
	#10 fw_in = 64'h0026_0024_002f_0012;
	#10 fw_in = 64'h004a_002c_0036_005c;


	#10 fw_in = 64'h0057_004f_005c_0045;
	#10 fw_in = 64'h0031_0029_001c_0014;
	#10 fw_in = 64'h0019_000c_005b_0019;
	#10 fw_in = 64'h0044_002c_0032_0003;
	#10 fw_in = 64'h0020_0026_000d_003a;
	#10 fw_in = 64'h0033_0000_005c_0051;
	#10 fw_in = 64'h0050_0063_0031_0023;
	#10 fw_in = 64'h001d_000b_0028_0060;


	#10 fw_in = 64'h000b_005c_001a_001d;
	#10 fw_in = 64'h0040_0025_0012_0013;
	#10 fw_in = 64'h001f_003b_005b_0038;
	#10 fw_in = 64'h0022_003e_0048_0005;
	#10 fw_in = 64'h0005_004a_005a_0056;
	#10 fw_in = 64'h0000_0033_0006_0034;
	#10 fw_in = 64'h0007_0056_0004_0045;
	#10 fw_in = 64'h0015_0032_0028_0060;


	#10 fw_in = 64'h002a_0059_0051_0044;
	#10 fw_in = 64'h000c_0005_0042_0047;
	#10 fw_in = 64'h005b_0029_0055_0001;
	#10 fw_in = 64'h0059_0028_005b_0003;
	#10 fw_in = 64'h003f_005a_0050_000f;
	#10 fw_in = 64'h0000_005f_004c_0013;
	#10 fw_in = 64'h005b_0010_0018_0029;
	#10 fw_in = 64'h0009_001d_001a_0064;


	#10 fw_in = 64'h004e_0040_001b_0044;
	#10 fw_in = 64'h003d_0042_0052_0061;
	#10 fw_in = 64'h0013_0047_0038_0025;
	#10 fw_in = 64'h0061_0021_002b_000c;
	#10 fw_in = 64'h0055_0047_0016_0050;
	#10 fw_in = 64'h0029_0023_001c_0049;
	#10 fw_in = 64'h0063_0049_0054_0000;
	#10 fw_in = 64'h0033_0030_0040_001f;


	#10 fw_in = 64'h0042_0055_0039_001e;
	#10 fw_in = 64'h0017_0013_003c_0045;
	#10 fw_in = 64'h000a_0044_004d_0025;
	#10 fw_in = 64'h005d_0003_0004_0007;
	#10 fw_in = 64'h0053_0054_000b_0045;
	#10 fw_in = 64'h0045_0012_0038_0016;
	#10 fw_in = 64'h0037_0035_0019_0000;
	#10 fw_in = 64'h005e_0028_005b_003f;


	#10 fw_in = 64'h003c_000f_004a_001f;
	#10 fw_in = 64'h0053_0019_0030_0017;
	#10 fw_in = 64'h0037_0005_0021_0024;
	#10 fw_in = 64'h0029_0057_0063_002c;
	#10 fw_in = 64'h003f_003f_003c_004f;
	#10 fw_in = 64'h0018_0031_002a_0054;
	#10 fw_in = 64'h0017_0049_0000_0019;
	#10 fw_in = 64'h003a_0016_0024_0037;


	#10 fw_in = 64'h005a_0004_004a_0053;
	#10 fw_in = 64'h001d_001d_0025_0009;
	#10 fw_in = 64'h0052_0006_002b_0035;
	#10 fw_in = 64'h0060_001d_0022_0055;
	#10 fw_in = 64'h005b_0008_0046_0006;
	#10 fw_in = 64'h0004_002f_000f_0047;
	#10 fw_in = 64'h0033_0048_0000_0054;
	#10 fw_in = 64'h004f_0063_0025_0062;


	#10 fw_in = 64'h004d_0048_0030_0042;
	#10 fw_in = 64'h0004_0002_0013_0046;
	#10 fw_in = 64'h003c_0008_0022_0036;
	#10 fw_in = 64'h0015_0062_0007_001d;
	#10 fw_in = 64'h0063_0023_0009_0055;
	#10 fw_in = 64'h0010_0063_004d_005c;
	#10 fw_in = 64'h005a_0000_0048_0035;
	#10 fw_in = 64'h0011_000b_0007_003c;


	#10 fw_in = 64'h002d_0034_003f_001f;
	#10 fw_in = 64'h0064_0059_0021_0010;
	#10 fw_in = 64'h0014_001d_0025_0064;
	#10 fw_in = 64'h002c_0004_0040_0016;
	#10 fw_in = 64'h005d_004f_005a_003b;
	#10 fw_in = 64'h0056_0024_005a_003f;
	#10 fw_in = 64'h0020_0000_0049_0049;
	#10 fw_in = 64'h0062_0059_003d_0054;


	#10 fw_in = 64'h0001_0028_000a_0019;
	#10 fw_in = 64'h0052_0036_000a_004f;
	#10 fw_in = 64'h001b_005a_0027_000f;
	#10 fw_in = 64'h0058_0018_0030_0044;
	#10 fw_in = 64'h0052_0017_0021_0020;
	#10 fw_in = 64'h005b_0050_0033_004c;
	#10 fw_in = 64'h0000_0020_0033_0037;
	#10 fw_in = 64'h0052_005f_003a_000e;


	#10 fw_in = 64'h0014_0037_0047_003f;
	#10 fw_in = 64'h002c_0046_0034_0029;
	#10 fw_in = 64'h0025_001c_0008_0050;
	#10 fw_in = 64'h002d_0001_0062_002b;
	#10 fw_in = 64'h005c_003a_004b_000d;
	#10 fw_in = 64'h0007_0026_0045_000d;
	#10 fw_in = 64'h0000_005a_0017_0063;
	#10 fw_in = 64'h0038_000b_0013_004d;


	#10 fw_in = 64'h0022_0015_0004_0052;
	#10 fw_in = 64'h0010_0058_0052_0053;
	#10 fw_in = 64'h0017_0005_001a_0061;
	#10 fw_in = 64'h0021_0062_0034_005d;
	#10 fw_in = 64'h0010_0007_0052_0023;
	#10 fw_in = 64'h0064_0060_0009_003a;
	#10 fw_in = 64'h004d_0054_0062_003f;
	#10 fw_in = 64'h000a_004e_0037_0000;


	#10 fw_in = 64'h0029_0064_0061_0018;
	#10 fw_in = 64'h002f_0012_0026_0032;
	#10 fw_in = 64'h0021_0033_002e_0033;
	#10 fw_in = 64'h001e_0052_0036_0045;
	#10 fw_in = 64'h003a_000f_0038_0057;
	#10 fw_in = 64'h0060_005c_005e_0050;
	#10 fw_in = 64'h000e_003c_0037_001f;
	#10 fw_in = 64'h0049_005e_002c_0000;


	#10 fw_in = 64'h0016_0053_0021_0058;
	#10 fw_in = 64'h0053_003d_0040_0043;
	#10 fw_in = 64'h0056_0057_0056_000c;
	#10 fw_in = 64'h000f_0054_005b_001f;
	#10 fw_in = 64'h005d_0015_0011_004d;
	#10 fw_in = 64'h001a_0028_001d_001a;
	#10 fw_in = 64'h0013_003d_0025_005b;
	#10 fw_in = 64'h001d_0026_0000_002c;


	#10 fw_in = 64'h001e_0021_0052_0044;
	#10 fw_in = 64'h0045_0012_001d_0061;
	#10 fw_in = 64'h0038_0055_0039_0045;
	#10 fw_in = 64'h005b_0030_005d_001d;
	#10 fw_in = 64'h0010_0048_002a_0001;
	#10 fw_in = 64'h0028_0036_0013_004e;
	#10 fw_in = 64'h003a_0007_0024_0040;
	#10 fw_in = 64'h004b_004e_0000_0037;


	#10 fw_in = 64'h0038_000b_0016_0053;
	#10 fw_in = 64'h0047_0010_001a_0059;
	#10 fw_in = 64'h0017_0009_0036_0026;
	#10 fw_in = 64'h0062_003a_0033_0054;
	#10 fw_in = 64'h0048_0046_001b_001c;
	#10 fw_in = 64'h001d_000b_0032_0034;
	#10 fw_in = 64'h000b_0059_0063_0028;
	#10 fw_in = 64'h005b_0000_004e_005e;


	#10 fw_in = 64'h0020_003d_0006_0024;
	#10 fw_in = 64'h0029_0061_004c_0018;
	#10 fw_in = 64'h005f_003b_0050_0048;
	#10 fw_in = 64'h0053_0027_0057_005a;
	#10 fw_in = 64'h0016_001e_0015_002f;
	#10 fw_in = 64'h0032_002c_0006_0056;
	#10 fw_in = 64'h005f_000b_0016_0030;
	#10 fw_in = 64'h002e_0000_0026_004e;


	#10 fw_in = 64'h0020_0035_0064_004d;
	#10 fw_in = 64'h003a_0064_004e_0058;
	#10 fw_in = 64'h002a_0012_0035_0043;
	#10 fw_in = 64'h0055_0063_0045_0024;
	#10 fw_in = 64'h0043_0006_004d_0060;
	#10 fw_in = 64'h0009_001d_0037_001d;
	#10 fw_in = 64'h0038_0062_004f_005e;
	#10 fw_in = 64'h0000_002e_004b_0049;


	#10 fw_in = 64'h0012_004d_001a_001e;
	#10 fw_in = 64'h0017_0019_0008_0013;
	#10 fw_in = 64'h0005_0015_0013_004a;
	#10 fw_in = 64'h0029_003c_001a_0049;
	#10 fw_in = 64'h003a_0001_0022_001b;
	#10 fw_in = 64'h0015_004a_0053_0025;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 0;
	#10 in_valid = 1;
	fw_in = 64'h0052_0011_003a_0033;
	#10 fw_in = 64'h0000_005b_001d_000a;

	#10 in_valid = 0;
end
endmodule
